library ieee;
use ieee.std_logic_1164.all; 
use ieee.std_logic_unsigned.all;

entity ROM_176x4 is
  port (Clock : in std_logic;
  		CS_L : in std_logic;
        R_W  : in std_logic;
        Addr   : in std_logic_vector(7 downto 0);
        Data  : out std_logic_vector(3 downto 0));
end ROM_176x4;

architecture ROM_176x4_Arch of ROM_176x4 is
  type rom_type is array (0 to 175)
        of std_logic_vector (3 downto 0);
  signal ROM : rom_type;
  signal Read_Enable : std_logic;
begin

ROM(0) <= X"7";
ROM(1) <= X"0";
ROM(2) <= X"D";
ROM(3) <= X"0";
ROM(4) <= X"B";
ROM(5) <= X"7";
ROM(6) <= X"9";
ROM(7) <= X"D";
ROM(8) <= X"1";
ROM(9) <= X"B";
ROM(10) <= X"0";
ROM(11) <= X"0";
ROM(12) <= X"0";
ROM(13) <= X"F";
ROM(14) <= X"0";
ROM(15) <= X"B";
ROM(16) <= X"4";
ROM(17) <= X"2";
ROM(18) <= X"F";
ROM(19) <= X"1";
ROM(20) <= X"B";
ROM(21) <= X"4";
ROM(22) <= X"1";
ROM(23) <= X"0";
ROM(24) <= X"5";
ROM(25) <= X"0";
ROM(26) <= X"B";
ROM(27) <= X"D";
ROM(28) <= X"4";
ROM(29) <= X"9";
ROM(30) <= X"3";
ROM(31) <= X"2";
ROM(32) <= X"0";
ROM(33) <= X"0";
ROM(34) <= X"0";
ROM(35) <= X"F";
ROM(36) <= X"0";
ROM(37) <= X"B";
ROM(38) <= X"6";
ROM(39) <= X"1";
ROM(40) <= X"D";
ROM(41) <= X"0";
ROM(42) <= X"B";
ROM(43) <= X"6";
ROM(44) <= X"6";
ROM(45) <= X"A";
ROM(46) <= X"5";
ROM(47) <= X"3";
ROM(48) <= X"9";
ROM(49) <= X"D";
ROM(50) <= X"0";
ROM(51) <= X"0";
ROM(52) <= X"0";
ROM(53) <= X"7";
ROM(54) <= X"0";
ROM(55) <= X"D";
ROM(56) <= X"0";
ROM(57) <= X"B";
ROM(58) <= X"F";
ROM(59) <= X"1";
ROM(60) <= X"B";
ROM(61) <= X"6";
ROM(62) <= X"1";
ROM(63) <= X"D";
ROM(64) <= X"1";
ROM(65) <= X"B";
ROM(66) <= X"6";
ROM(67) <= X"6";
ROM(68) <= X"A";
ROM(69) <= X"4";
ROM(70) <= X"7";
ROM(71) <= X"9";
ROM(72) <= X"D";
ROM(73) <= X"0";
ROM(74) <= X"0";
ROM(75) <= X"0";
ROM(76) <= X"0";
ROM(77) <= X"F";
ROM(78) <= X"0";
ROM(79) <= X"B";
ROM(80) <= X"6";
ROM(81) <= X"F";
ROM(82) <= X"D";
ROM(83) <= X"0";
ROM(84) <= X"B";
ROM(85) <= X"A";
ROM(86) <= X"C";
ROM(87) <= X"5";
ROM(88) <= X"9";
ROM(89) <= X"D";
ROM(90) <= X"0";
ROM(91) <= X"0";
ROM(92) <= X"4";
ROM(93) <= X"2";
ROM(94) <= X"7";
ROM(95) <= X"9";
ROM(96) <= X"D";
ROM(97) <= X"0";
ROM(98) <= X"B";
ROM(99) <= X"F";
ROM(100) <= X"1";
ROM(101) <= X"B";
ROM(102) <= X"6";
ROM(103) <= X"F";
ROM(104) <= X"D";
ROM(105) <= X"1";
ROM(106) <= X"B";
ROM(107) <= X"6";
ROM(108) <= X"1";
ROM(109) <= X"A";
ROM(110) <= X"F";
ROM(111) <= X"7";
ROM(112) <= X"9";
ROM(113) <= X"D";
ROM(114) <= X"0";
ROM(115) <= X"0";
ROM(116) <= X"7";
ROM(117) <= X"0";
ROM(118) <= X"D";
ROM(119) <= X"0";
ROM(120) <= X"B";
ROM(121) <= X"D";
ROM(122) <= X"1";
ROM(123) <= X"B";
ROM(124) <= X"9";
ROM(125) <= X"D";
ROM(126) <= X"0";
ROM(127) <= X"7";
ROM(128) <= X"9";
ROM(129) <= X"D";
ROM(130) <= X"0";
ROM(131) <= X"B";
ROM(132) <= X"D";
ROM(133) <= X"1";
ROM(134) <= X"B";
ROM(135) <= X"9";
ROM(136) <= X"D";
ROM(137) <= X"0";
ROM(138) <= X"0";
ROM(139) <= X"0";
ROM(140) <= X"0";
ROM(141) <= X"0";
ROM(142) <= X"0";
ROM(143) <= X"0";
ROM(144) <= X"0";
ROM(145) <= X"0";
ROM(146) <= X"0";
ROM(147) <= X"0";
ROM(148) <= X"0";
ROM(149) <= X"0";
ROM(150) <= X"0";
ROM(151) <= X"0";
ROM(152) <= X"0";
ROM(153) <= X"0";
ROM(154) <= X"0";
ROM(155) <= X"0";
ROM(156) <= X"0";
ROM(157) <= X"0";
ROM(158) <= X"0";
ROM(159) <= X"0";
ROM(160) <= X"0";
ROM(161) <= X"0";
ROM(162) <= X"0";
ROM(163) <= X"0";
ROM(164) <= X"0";
ROM(165) <= X"0";
ROM(166) <= X"0";
ROM(167) <= X"0";
ROM(168) <= X"0";
ROM(169) <= X"0";
ROM(170) <= X"0";
ROM(171) <= X"0";
ROM(172) <= X"0";
ROM(173) <= X"0";
ROM(174) <= X"0";
ROM(175) <= X"0";
	Read_Enable <=  '0' when(CS_L='0' and R_W = '1') else '1';

	process (Clock)
	begin
		if(Clock='0') then
			if(Read_Enable = '0') then
			  Data  <= ROM(conv_integer(Addr));
		  	else
			  Data <= "ZZZZ";
	      	end if;
		else Data <= "ZZZZ";
		end if;

	end process;

	end ROM_176x4_Arch;
